module foo();
   reg

endmodule
