module module4 (
    input wire a,
    output wire b
);

    assign b = ~a;

endmodule
